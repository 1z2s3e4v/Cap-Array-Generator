* SPICE NETLIST
***************************************

.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT cfmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_wo PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_2t PLUS MINUS
.ENDS
***************************************
.SUBCKT cfmom_mx_4t PLUS1 MINUS1 PLUS2 MINUS2
.ENDS
***************************************
.SUBCKT cfmom_wo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT cfmom_wo_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT cmoscap_rf GATE BULK GNODE
.ENDS
***************************************
.SUBCKT cmoscap_rf18 GATE BULK GNODE
.ENDS
***************************************
.SUBCKT cmoscap_rf18_nw GATE BULK GNODE
.ENDS
***************************************
.SUBCKT cmoscap_rf25 GATE BULK GNODE
.ENDS
***************************************
.SUBCKT cmoscap_rf25_nw GATE BULK GNODE
.ENDS
***************************************
.SUBCKT cmoscap_rf_nw GATE BULK GNODE
.ENDS
***************************************
.SUBCKT dmoscap_rf GATE1 GATE2 BULK GNODE
.ENDS
***************************************
.SUBCKT dmoscap_rf18 GATE1 GATE2 BULK GNODE
.ENDS
***************************************
.SUBCKT dmoscap_rf18_nw GATE1 GATE2 BULK GNODE
.ENDS
***************************************
.SUBCKT dmoscap_rf25 GATE1 GATE2 BULK GNODE
.ENDS
***************************************
.SUBCKT dmoscap_rf25_nw GATE1 GATE2 BULK GNODE
.ENDS
***************************************
.SUBCKT dmoscap_rf_nw GATE1 GATE2 BULK GNODE
.ENDS
***************************************
.SUBCKT mimcap_sin TOP BOTTOM
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf15_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ndio_gated_mac PLUS MINUS
.ENDS
***************************************
.SUBCKT ndio_hia_mac PLUS MINUS
.ENDS
***************************************
.SUBCKT ndio_hia_rf CATHODE ANODE
.ENDS
***************************************
.SUBCKT nmos_rf_18_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18ud15_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_18ud15_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18ud15_nw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_25_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_nw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_nw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_ulvt_5t D G S B NG
.ENDS
***************************************
.SUBCKT nmos_rf_ulvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_ulvt_nw D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_15 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_edc PLUS MINUS
.ENDS
***************************************
.SUBCKT pcmoscap_rf GATE BULK GNODE
.ENDS
***************************************
.SUBCKT pcmoscap_rf18 GATE BULK GNODE
.ENDS
***************************************
.SUBCKT pcmoscap_rf25 GATE BULK GNODE
.ENDS
***************************************
.SUBCKT pdio_gated_mac PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_gated_mac_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pdio_hia_mac PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_hia_rf ANODE CATHODE GNODE
.ENDS
***************************************
.SUBCKT pmos_rf_18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18ud15_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18ud15_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18ud15_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_ulvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_ulvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_ulvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT pmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmoscap_rf GATE BULK GNODE
.ENDS
***************************************
.SUBCKT pmoscap_rf18 GATE BULK GNODE
.ENDS
***************************************
.SUBCKT probe1 TOP BULK
.ENDS
***************************************
.SUBCKT probe2 TOP BULK
.ENDS
***************************************
.SUBCKT probe3 TOP BULK
.ENDS
***************************************
.SUBCKT probe4 TOP BULK
.ENDS
***************************************
.SUBCKT probe5 TOP BULK
.ENDS
***************************************
.SUBCKT probe6 TOP BULK
.ENDS
***************************************
.SUBCKT probe7 TOP BULK
.ENDS
***************************************
.SUBCKT rm1w PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2w PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3w PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4w PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5w PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6w PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7w PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8w PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9w PLUS MINUS
.ENDS
***************************************
.SUBCKT rmap PLUS MINUS
.ENDS
***************************************
.SUBCKT rnmg PLUS MINUS
.ENDS
***************************************
.SUBCKT rnmg_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpmg PLUS MINUS
.ENDS
***************************************
.SUBCKT rpmg_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rupolym PLUS MINUS
.ENDS
***************************************
.SUBCKT rupolym_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rupolym_rf HI LO GNODE
.ENDS
***************************************
.SUBCKT spiral_std_mu_a28_dm TOP BOTTOM GNODE
.ENDS
***************************************
.SUBCKT spiral_std_mu_z TOP BOTTOM GNODE
.ENDS
***************************************
.SUBCKT spiral_std_mu_z_dm TOP BOTTOM GNODE
.ENDS
***************************************
.SUBCKT spiral_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_lc PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_a28_a28_dm TOP BOTTOM GNODE TAP
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z_a TOP BOTTOM GNODE TAP
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z_a28_dm TOP BOTTOM GNODE TAP
.ENDS
***************************************
.SUBCKT spiral_sym_ct_rl PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_a28_dm TOP BOTTOM GNODE
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z TOP BOTTOM GNODE
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z_dm TOP BOTTOM GNODE
.ENDS
***************************************
.SUBCKT CU1F 1 2
** N=4 EP=2 IP=0 FDC=1
X0 2 1 cfmom_2t w=1.2e-06 s=5e-08 nr=3 lr=2.29417e-06 stm=4 spm=6 $X=0 $Y=2100 $D=656
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3
** N=5 EP=3 IP=8 FDC=2
X0 1 2 CU1F $T=0 0 0 0 $X=-350 $Y=0
X1 3 2 CU1F $T=2100 0 0 0 $X=1750 $Y=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5
** N=7 EP=5 IP=10 FDC=4
X0 1 3 2 ICV_1 $T=0 0 0 0 $X=-350 $Y=0
X1 4 3 5 ICV_1 $T=4200 0 0 0 $X=3850 $Y=0
.ENDS
***************************************
.SUBCKT ARRAY_CMP_T1 SL3A SL3B SL2A SL2B SL1A SL1B VSS09A TOP_ARRAY VDD09A
** N=11 EP=9 IP=46 FDC=22
X0 VSS09A TOP_ARRAY CU1F $T=37800 0 0 0 $X=37450 $Y=0
X1 VDD09A VDD09A CU1F $T=45200 0 0 0 $X=44850 $Y=0
X2 SL3A TOP_ARRAY SL3A ICV_1 $T=33600 0 0 0 $X=33250 $Y=0
X3 VDD09A VDD09A VDD09A ICV_1 $T=41000 0 0 0 $X=40650 $Y=0
X4 VSS09A VSS09A TOP_ARRAY VSS09A VSS09A ICV_2 $T=0 0 0 0 $X=-350 $Y=0
X5 SL3A SL3A TOP_ARRAY SL3B SL3B ICV_2 $T=8400 0 0 0 $X=8050 $Y=0
X6 SL2A SL2B TOP_ARRAY SL1B SL1A ICV_2 $T=16800 0 0 0 $X=16450 $Y=0
X7 SL2B SL2A TOP_ARRAY SL3B SL3B ICV_2 $T=25200 0 0 0 $X=24850 $Y=0
.ENDS
***************************************
